../hw/vendor/esl_epfl_x_heep/tb/tb_util.svh